`timescale  1ns / 1ns
module INSTRUCTION_MEMORY (input [31:0] PC_out, output reg [31:0] INS_out);
  reg [31:0] mem [99:0];
  integer i;
  initial begin
    for(i=0; i<100; i=i+1) mem[i] = 32'b0;
    // INSERT INSTRUCTIONS HERE for example mem[0] = 000000 00011 00010 00001 00000 100000 (without spaces)
    // is for add $1, $2, $3

    mem[0]  = 32'b10001100000000010000001110000100;
    mem[1]  = 32'b10001100000000100000001110000101;
    mem[2]  = 32'b10001100000000110000001110000110;
    mem[3]  = 32'b10001100001001010000000000000000;
    mem[4]  = 32'b00010000001000100000000000001000;
    mem[5]  = 32'b00000000011000010000100000100000;
    mem[6]  = 32'b10001100001001000000000000000000;
    mem[7]  = 32'b00000000101001000011000000101010;
    mem[8]  = 32'b00000000000000000000000000000000;
    mem[9]  = 32'b00000000000000000000000000000000;
    mem[10]  = 32'b00010000000001100000000000000001;
    mem[11] = 32'b00000000000001000010100000100000;
    mem[12] = 32'b00001000000000000000000000000100;
  end

  always @ (PC_out) INS_out <= mem[PC_out];

endmodule
